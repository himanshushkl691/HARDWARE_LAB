module AND_32BIT(out,in0,in1);
   input[31:0] in0,in1;
   output [31:0] out;
   AND and0[31:0](out,in0,in1);
endmodule // AND_32BIT

