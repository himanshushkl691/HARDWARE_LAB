module ADDER_32BIT(sum,carry,a,b,cin);
   input[31:0] a,b;
   output [31:0] sum;
   input cin;
   output carry;
   FULL_ADDER fa1(sum[0],c,a[0],b[0],cin);
   FULL_ADDER fa2(sum[1],d,a[1],b[1],c);
   FULL_ADDER fa3(sum[2],e,a[2],b[2],d);
   FULL_ADDER fa4(sum[3],f,a[3],b[3],e);
   FULL_ADDER fa5(sum[4],g,a[4],b[4],f);
   FULL_ADDER fa6(sum[5],h,a[5],b[5],g);
   FULL_ADDER fa7(sum[6],i,a[6],b[6],h);
   FULL_ADDER fa8(sum[7],j,a[7],b[7],i);
   FULL_ADDER fa9(sum[8],k,a[8],b[8],j);
   FULL_ADDER fa10(sum[9],l,a[9],b[9],k);
   FULL_ADDER fa11(sum[10],m,a[10],b[10],l);
   FULL_ADDER fa12(sum[11],n,a[11],b[11],m);
   FULL_ADDER fa13(sum[12],o,a[12],b[12],n);
   FULL_ADDER fa14(sum[13],p,a[13],b[13],o);
   FULL_ADDER fa15(sum[14],q,a[14],b[14],p);
   FULL_ADDER fa16(sum[15],r,a[15],b[15],q);

   FULL_ADDER fa17(sum[16],s,a[16],b[16],r);
   FULL_ADDER fa18(sum[17],t,a[17],b[17],s);
   FULL_ADDER fa19(sum[18],u,a[18],b[18],t);
   FULL_ADDER fa20(sum[19],v,a[19],b[19],u);
   FULL_ADDER fa21(sum[20],w,a[20],b[20],v);
   FULL_ADDER fa22(sum[21],x,a[21],b[21],w);
   FULL_ADDER fa23(sum[22],y,a[22],b[22],x);
   FULL_ADDER fa24(sum[23],z,a[23],b[23],y);
   FULL_ADDER fa25(sum[24],a0,a[24],b[24],z);
   FULL_ADDER fa26(sum[25],b0,a[25],b[25],a0);
   FULL_ADDER fa27(sum[26],c0,a[26],b[26],b0);
   FULL_ADDER fa28(sum[27],d0,a[27],b[27],c0);
   FULL_ADDER fa29(sum[28],e0,a[28],b[28],d0);
   FULL_ADDER fa30(sum[29],f0,a[29],b[29],e0);
   FULL_ADDER fa31(sum[30],g0,a[30],b[30],f0);
   FULL_ADDER fa32(sum[31],carry,a[31],b[31],g0);
endmodule // ADDER_16BIT
